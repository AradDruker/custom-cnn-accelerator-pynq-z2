library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library xil_defaultlib;
use xil_defaultlib.types_package.all;

entity TB_layer_5 is
--  Port ( );
end TB_layer_5;

architecture Behavioral of TB_layer_5 is

	component layer_5 is
		Port (
			clka   : in  std_logic; -- Clock signal
			resetn : in  std_logic; -- Active-low reset signal
			start  : in  std_logic; -- Start signal to begin operation
			finish : out std_logic; -- Indicates when operation is complete

			bias : in bais_array(0 to 119); -- Bias to be added after convolution

			addrb_weights_fc1 : out address_array_weights_fc1(0 to 119);
			doutb_weights_fc1 : in  bram_data_array(0 to 119);

			--wea_layer_5   : out wea_array(0 to 11);
			--addra_layer_5 : out std_logic_vector(3 downto 0);
			--dina_layer_5  : out bram_data_array(0 to 11);

			wea_layer_5   : out std_logic_vector(0 downto 0);
			addra_layer_5 : out std_logic_vector(6 downto 0);
			dina_layer_5  : out std_logic_vector(7 downto 0);

			addrb_layer_4 : out address_array_layer_4(0 to 15);
			doutb_layer_4 : in  bram_data_array(0 to 15);
			locked_debug  : out std_logic
		);
	end component;

	signal clka         : std_logic := '0';
	signal resetn       : std_logic := '1';
	signal start        : std_logic := '0';
	signal finish       : std_logic;
	signal locked_debug : std_logic;

	signal bias : bais_array(0 to 119) := (others => to_signed(-40, 32));

	constant CLK_PERIOD : time := 10 ns;

	signal resetn_flag : integer := 0;
	signal start_flag  : integer := 0;

	signal wea_layer_5   : std_logic_vector(0 downto 0);
	signal addra_layer_5 : std_logic_vector(6 downto 0);
	signal dina_layer_5  : std_logic_vector(7 downto 0);

	signal addrb_layer_4     : address_array_layer_4(0 to 15);
	signal addrb_weights_fc1 : address_array_weights_fc1(0 to 119);
	signal doutb_layer_4     : bram_data_array(0 to 15);
	signal doutb_weights_fc1 : bram_data_array(0 to 119);

	signal inputs : bram_data_array(0 to 399) := (
			std_logic_vector(to_unsigned( 17 , 8)),
			std_logic_vector(to_unsigned( 31 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 21 , 8)),
			std_logic_vector(to_unsigned( 14 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 42 , 8)),
			std_logic_vector(to_unsigned( 59 , 8)),
			std_logic_vector(to_unsigned( 51 , 8)),
			std_logic_vector(to_unsigned( 12 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 63 , 8)),
			std_logic_vector(to_unsigned( 76 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 17 , 8)),
			std_logic_vector(to_unsigned( 44 , 8)),
			std_logic_vector(to_unsigned( 73 , 8)),
			std_logic_vector(to_unsigned( 26 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 12 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 19 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 7 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 23 , 8)),
			std_logic_vector(to_unsigned( 28 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 18 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 36 , 8)),
			std_logic_vector(to_unsigned( 40 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 29 , 8)),
			std_logic_vector(to_unsigned( 11 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 22 , 8)),
			std_logic_vector(to_unsigned( 13 , 8)),
			std_logic_vector(to_unsigned( 1 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 19 , 8)),
			std_logic_vector(to_unsigned( 19 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 56 , 8)),
			std_logic_vector(to_unsigned( 53 , 8)),
			std_logic_vector(to_unsigned( 44 , 8)),
			std_logic_vector(to_unsigned( 54 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 22 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 31 , 8)),
			std_logic_vector(to_unsigned( 51 , 8)),
			std_logic_vector(to_unsigned( 31 , 8)),
			std_logic_vector(to_unsigned( 23 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 18 , 8)),
			std_logic_vector(to_unsigned( 42 , 8)),
			std_logic_vector(to_unsigned( 18 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 40 , 8)),
			std_logic_vector(to_unsigned( 30 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 38 , 8)),
			std_logic_vector(to_unsigned( 26 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 35 , 8)),
			std_logic_vector(to_unsigned( 31 , 8)),
			std_logic_vector(to_unsigned( 41 , 8)),
			std_logic_vector(to_unsigned( 68 , 8)),
			std_logic_vector(to_unsigned( 37 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 19 , 8)),
			std_logic_vector(to_unsigned( 38 , 8)),
			std_logic_vector(to_unsigned( 14 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 30 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 20 , 8)),
			std_logic_vector(to_unsigned( 14 , 8)),
			std_logic_vector(to_unsigned( 13 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 20 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 5 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 7 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 20 , 8)),
			std_logic_vector(to_unsigned( 21 , 8)),
			std_logic_vector(to_unsigned( 17 , 8)),
			std_logic_vector(to_unsigned( 23 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 25 , 8)),
			std_logic_vector(to_unsigned( 33 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 64 , 8)),
			std_logic_vector(to_unsigned( 54 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 72 , 8)),
			std_logic_vector(to_unsigned( 49 , 8)),
			std_logic_vector(to_unsigned( 1 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 48 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 80 , 8)),
			std_logic_vector(to_unsigned( 115 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 44 , 8)),
			std_logic_vector(to_unsigned( 121 , 8)),
			std_logic_vector(to_unsigned( 86 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 120 , 8)),
			std_logic_vector(to_unsigned( 127 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 23 , 8)),
			std_logic_vector(to_unsigned( 106 , 8)),
			std_logic_vector(to_unsigned( 55 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 22 , 8)),
			std_logic_vector(to_unsigned( 41 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 5 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 43 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 5 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 50 , 8)),
			std_logic_vector(to_unsigned( 54 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 18 , 8)),
			std_logic_vector(to_unsigned( 9 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 11 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 4 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 26 , 8)),
			std_logic_vector(to_unsigned( 24 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 8 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 28 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 45 , 8)),
			std_logic_vector(to_unsigned( 37 , 8)),
			std_logic_vector(to_unsigned( 54 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 25 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 26 , 8)),
			std_logic_vector(to_unsigned( 31 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 5 , 8)),
			std_logic_vector(to_unsigned( 9 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 20 , 8)),
			std_logic_vector(to_unsigned( 2 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 24 , 8)),
			std_logic_vector(to_unsigned( 10 , 8)),
			std_logic_vector(to_unsigned( 12 , 8)),
			std_logic_vector(to_unsigned( 23 , 8)),
			std_logic_vector(to_unsigned( 32 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 35 , 8)),
			std_logic_vector(to_unsigned( 30 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 7 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 16 , 8)),
			std_logic_vector(to_unsigned( 36 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 21 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 1 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 15 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 13 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 3 , 8)),
			std_logic_vector(to_unsigned( 25 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 22 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 22 , 8)),
			std_logic_vector(to_unsigned( 7 , 8)),
			std_logic_vector(to_unsigned( 33 , 8)),
			std_logic_vector(to_unsigned( 86 , 8)),
			std_logic_vector(to_unsigned( 1 , 8)),
			std_logic_vector(to_unsigned( 9 , 8)),
			std_logic_vector(to_unsigned( 6 , 8)),
			std_logic_vector(to_unsigned( 75 , 8)),
			std_logic_vector(to_unsigned( 104 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 61 , 8)),
			std_logic_vector(to_unsigned( 53 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 38 , 8)),
			std_logic_vector(to_unsigned( 58 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 34 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8)),
			std_logic_vector(to_unsigned( 0 , 8))
	);
	signal weights : bram_data_array(0 to 399) := (
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 32 , 8)),
			std_logic_vector(to_signed( 36 , 8)),
			std_logic_vector(to_signed( 30 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( -29 , 8)),
			std_logic_vector(to_signed( 11 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( -20 , 8)),
			std_logic_vector(to_signed( -9 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( -25 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 27 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( -40 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( -25 , 8)),
			std_logic_vector(to_signed( -45 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( 38 , 8)),
			std_logic_vector(to_signed( 41 , 8)),
			std_logic_vector(to_signed( 43 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 28 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 20 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 28 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( 21 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -32 , 8)),
			std_logic_vector(to_signed( -12 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 25 , 8)),
			std_logic_vector(to_signed( 32 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( -48 , 8)),
			std_logic_vector(to_signed( -32 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( 46 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( -20 , 8)),
			std_logic_vector(to_signed( 16 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( -28 , 8)),
			std_logic_vector(to_signed( -17 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( -12 , 8)),
			std_logic_vector(to_signed( -47 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 30 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( 33 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( -21 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( -14 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( -26 , 8)),
			std_logic_vector(to_signed( -9 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -24 , 8)),
			std_logic_vector(to_signed( -25 , 8)),
			std_logic_vector(to_signed( -19 , 8)),
			std_logic_vector(to_signed( 16 , 8)),
			std_logic_vector(to_signed( 16 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( -19 , 8)),
			std_logic_vector(to_signed( 31 , 8)),
			std_logic_vector(to_signed( 23 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( -15 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( -27 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -15 , 8)),
			std_logic_vector(to_signed( -12 , 8)),
			std_logic_vector(to_signed( -15 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -33 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( -18 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 27 , 8)),
			std_logic_vector(to_signed( 30 , 8)),
			std_logic_vector(to_signed( 27 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 29 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 16 , 8)),
			std_logic_vector(to_signed( -50 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( -27 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( 10 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( -35 , 8)),
			std_logic_vector(to_signed( -35 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( -67 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 22 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( -27 , 8)),
			std_logic_vector(to_signed( -12 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 24 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( -42 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( -19 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( -18 , 8)),
			std_logic_vector(to_signed( -34 , 8)),
			std_logic_vector(to_signed( -29 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( -18 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 10 , 8)),
			std_logic_vector(to_signed( -23 , 8)),
			std_logic_vector(to_signed( -36 , 8)),
			std_logic_vector(to_signed( -21 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( -41 , 8)),
			std_logic_vector(to_signed( 11 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( -12 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 11 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( -6 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( -26 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -14 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( 21 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( 25 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 2 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( -14 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( 21 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( -21 , 8)),
			std_logic_vector(to_signed( -29 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( 3 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( -28 , 8)),
			std_logic_vector(to_signed( -19 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 26 , 8)),
			std_logic_vector(to_signed( -31 , 8)),
			std_logic_vector(to_signed( -49 , 8)),
			std_logic_vector(to_signed( -41 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 25 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( -27 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( -41 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( 20 , 8)),
			std_logic_vector(to_signed( 29 , 8)),
			std_logic_vector(to_signed( -19 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -14 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( 27 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( 12 , 8)),
			std_logic_vector(to_signed( 9 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( 29 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 29 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( 5 , 8)),
			std_logic_vector(to_signed( -15 , 8)),
			std_logic_vector(to_signed( -24 , 8)),
			std_logic_vector(to_signed( -16 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( 8 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 10 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( -8 , 8)),
			std_logic_vector(to_signed( -26 , 8)),
			std_logic_vector(to_signed( 15 , 8)),
			std_logic_vector(to_signed( 28 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( 22 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -11 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -13 , 8)),
			std_logic_vector(to_signed( -2 , 8)),
			std_logic_vector(to_signed( -9 , 8)),
			std_logic_vector(to_signed( -4 , 8)),
			std_logic_vector(to_signed( -17 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -14 , 8)),
			std_logic_vector(to_signed( -10 , 8)),
			std_logic_vector(to_signed( 6 , 8)),
			std_logic_vector(to_signed( -15 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( 14 , 8)),
			std_logic_vector(to_signed( 24 , 8)),
			std_logic_vector(to_signed( 32 , 8)),
			std_logic_vector(to_signed( 13 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( 0 , 8)),
			std_logic_vector(to_signed( 18 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( -42 , 8)),
			std_logic_vector(to_signed( 1 , 8)),
			std_logic_vector(to_signed( -3 , 8)),
			std_logic_vector(to_signed( -17 , 8)),
			std_logic_vector(to_signed( 19 , 8)),
			std_logic_vector(to_signed( -7 , 8)),
			std_logic_vector(to_signed( 17 , 8)),
			std_logic_vector(to_signed( -5 , 8)),
			std_logic_vector(to_signed( 7 , 8)),
			std_logic_vector(to_signed( 27 , 8)),
			std_logic_vector(to_signed( -34 , 8)),
			std_logic_vector(to_signed( 4 , 8)),
			std_logic_vector(to_signed( 11 , 8)),
			std_logic_vector(to_signed( -1 , 8)),
			std_logic_vector(to_signed( -22 , 8)),
			std_logic_vector(to_signed( -17 , 8))
	);

begin

		U1 : layer_5 port map(
			clka              => clka,
			resetn            => resetn,
			start             => start,
			finish            => finish,
			bias              => bias,
			addrb_weights_fc1 => addrb_weights_fc1,
			doutb_weights_fc1 => doutb_weights_fc1,
			wea_layer_5       => wea_layer_5,
			addra_layer_5     => addra_layer_5,
			dina_layer_5      => dina_layer_5,
			addrb_layer_4     => addrb_layer_4,
			doutb_layer_4     => doutb_layer_4,
			locked_debug      => locked_debug
		);

	clka_process : process
	begin
		while true loop
			clka <= '0';
			wait for CLK_PERIOD / 2;
			clka <= '1';
			wait for CLK_PERIOD / 2;
		end loop;
	end process;

	resetn_process : process(clka)
	begin
		if rising_edge(clka) then
			if resetn_flag = 0 then
				resetn      <= '0';
				resetn_flag <= 1;
			else
				resetn <= '1';
			end if;
		end if;
	end process;

	start_process : process(clka)
	begin
		if rising_edge(clka) and resetn = '1' then
			if start_flag = 0 and locked_debug = '1' then
				start      <= '1';
				start_flag <= 1;
			else
				start <= '0';
			end if;
		end if;
	end process;

	main_process : process(clka)
		variable index_weights : integer;
		variable index_inputs  : integer;
		variable bram_counter  : integer := 0;

	begin
		if resetn = '1' then
			if rising_edge(clka) then
				index_weights := to_integer(unsigned(addrb_weights_fc1(0)));

				if index_inputs = 24 and bram_counter < 15 then
					bram_counter := bram_counter + 1;
				end if;

				index_inputs := to_integer(unsigned(addrb_layer_4(bram_counter)));

				for i in 0 to 119 loop
					doutb_weights_fc1(i) <= weights(index_weights);
				end loop;

				doutb_layer_4(0)  <= inputs(index_inputs);
				doutb_layer_4(1)  <= inputs(1*25 + index_inputs);
				doutb_layer_4(2)  <= inputs(2*25 + index_inputs);
				doutb_layer_4(3)  <= inputs(3*25 + index_inputs);
				doutb_layer_4(4)  <= inputs(4*25 + index_inputs);
				doutb_layer_4(5)  <= inputs(5*25 + index_inputs);
				doutb_layer_4(6)  <= inputs(6*25 + index_inputs);
				doutb_layer_4(7)  <= inputs(7*25 + index_inputs);
				doutb_layer_4(8)  <= inputs(8*25 + index_inputs);
				doutb_layer_4(9)  <= inputs(9*25 + index_inputs);
				doutb_layer_4(10) <= inputs(10*25 + index_inputs);
				doutb_layer_4(11) <= inputs(11*25 + index_inputs);
				doutb_layer_4(12) <= inputs(12*25 + index_inputs);
				doutb_layer_4(13) <= inputs(13*25 + index_inputs);
				doutb_layer_4(14) <= inputs(14*25 + index_inputs);
				doutb_layer_4(15) <= inputs(15*25 + index_inputs);

			end if;
		end if;
	end process;

end Behavioral;