library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

library xil_defaultlib;
use xil_defaultlib.types_package.all;

entity TB_channel_layer_5 is
--  Port ( );
end TB_channel_layer_5;

architecture Behavioral of TB_channel_layer_5 is

	component channel_layer_5 is
		Port (
			clka   : in  std_logic; -- Clock signal
			resetn : in  std_logic; -- Active-low reset signal
			start  : in  std_logic; -- Start signal to begin operation
			finish : out std_logic; -- Indicates when operation is complete

			weight : in signed(7 downto 0);  -- Kernel weights for convolution
			bias   : in signed(31 downto 0); -- Bias to be added after convolution

			compute_output : out std_logic_vector(7 downto 0);
			data           : in  unsigned(7 downto 0);
			scale          : in  integer
		);
	end component;

	signal clka   : std_logic := '0';
	signal resetn : std_logic := '1';
	signal start  : std_logic := '0';
	signal finish : std_logic;

	constant CLK_PERIOD : time := 10 ns;

	signal resetn_flag    : integer := 0;
	signal start_flag     : integer := 0;
	signal compute_output : std_logic_vector(7 downto 0);

	signal weights : kernel_array(0 to 399) := (
			to_signed( 14 , 8),
			to_signed( -31 , 8),
			to_signed( -29 , 8),
			to_signed( -22 , 8),
			to_signed( -11 , 8),
			to_signed( 7 , 8),
			to_signed( -3 , 8),
			to_signed( 2 , 8),
			to_signed( -12 , 8),
			to_signed( -21 , 8),
			to_signed( 11 , 8),
			to_signed( 14 , 8),
			to_signed( 16 , 8),
			to_signed( 6 , 8),
			to_signed( 11 , 8),
			to_signed( -2 , 8),
			to_signed( -3 , 8),
			to_signed( 3 , 8),
			to_signed( 16 , 8),
			to_signed( 17 , 8),
			to_signed( 11 , 8),
			to_signed( -1 , 8),
			to_signed( -24 , 8),
			to_signed( 12 , 8),
			to_signed( 32 , 8),
			to_signed( -24 , 8),
			to_signed( 21 , 8),
			to_signed( 33 , 8),
			to_signed( 19 , 8),
			to_signed( 54 , 8),
			to_signed( -51 , 8),
			to_signed( -13 , 8),
			to_signed( -10 , 8),
			to_signed( 13 , 8),
			to_signed( 22 , 8),
			to_signed( -20 , 8),
			to_signed( -5 , 8),
			to_signed( -30 , 8),
			to_signed( -27 , 8),
			to_signed( -13 , 8),
			to_signed( -33 , 8),
			to_signed( 2 , 8),
			to_signed( 3 , 8),
			to_signed( 10 , 8),
			to_signed( -28 , 8),
			to_signed( -37 , 8),
			to_signed( 18 , 8),
			to_signed( 27 , 8),
			to_signed( 5 , 8),
			to_signed( -8 , 8),
			to_signed( 17 , 8),
			to_signed( 6 , 8),
			to_signed( 33 , 8),
			to_signed( 4 , 8),
			to_signed( 9 , 8),
			to_signed( 3 , 8),
			to_signed( 17 , 8),
			to_signed( 29 , 8),
			to_signed( 14 , 8),
			to_signed( 9 , 8),
			to_signed( -8 , 8),
			to_signed( 22 , 8),
			to_signed( 2 , 8),
			to_signed( 21 , 8),
			to_signed( 10 , 8),
			to_signed( -29 , 8),
			to_signed( 21 , 8),
			to_signed( 31 , 8),
			to_signed( 47 , 8),
			to_signed( -3 , 8),
			to_signed( -48 , 8),
			to_signed( -42 , 8),
			to_signed( -42 , 8),
			to_signed( -28 , 8),
			to_signed( -13 , 8),
			to_signed( 3 , 8),
			to_signed( -23 , 8),
			to_signed( -13 , 8),
			to_signed( -31 , 8),
			to_signed( -6 , 8),
			to_signed( 31 , 8),
			to_signed( 27 , 8),
			to_signed( 10 , 8),
			to_signed( 4 , 8),
			to_signed( -14 , 8),
			to_signed( 16 , 8),
			to_signed( 17 , 8),
			to_signed( 8 , 8),
			to_signed( 0 , 8),
			to_signed( -10 , 8),
			to_signed( 37 , 8),
			to_signed( 14 , 8),
			to_signed( 2 , 8),
			to_signed( -23 , 8),
			to_signed( -38 , 8),
			to_signed( -1 , 8),
			to_signed( 11 , 8),
			to_signed( 19 , 8),
			to_signed( -3 , 8),
			to_signed( -9 , 8),
			to_signed( -27 , 8),
			to_signed( -14 , 8),
			to_signed( 3 , 8),
			to_signed( -4 , 8),
			to_signed( -1 , 8),
			to_signed( 27 , 8),
			to_signed( 31 , 8),
			to_signed( 4 , 8),
			to_signed( -1 , 8),
			to_signed( -15 , 8),
			to_signed( -18 , 8),
			to_signed( 13 , 8),
			to_signed( 23 , 8),
			to_signed( 15 , 8),
			to_signed( 14 , 8),
			to_signed( -19 , 8),
			to_signed( -7 , 8),
			to_signed( -9 , 8),
			to_signed( -3 , 8),
			to_signed( -52 , 8),
			to_signed( -62 , 8),
			to_signed( -10 , 8),
			to_signed( -1 , 8),
			to_signed( -39 , 8),
			to_signed( -26 , 8),
			to_signed( -25 , 8),
			to_signed( -19 , 8),
			to_signed( -11 , 8),
			to_signed( -7 , 8),
			to_signed( 36 , 8),
			to_signed( -18 , 8),
			to_signed( -9 , 8),
			to_signed( -5 , 8),
			to_signed( -19 , 8),
			to_signed( -5 , 8),
			to_signed( 16 , 8),
			to_signed( 2 , 8),
			to_signed( 31 , 8),
			to_signed( 6 , 8),
			to_signed( -14 , 8),
			to_signed( -28 , 8),
			to_signed( 0 , 8),
			to_signed( -3 , 8),
			to_signed( -30 , 8),
			to_signed( -53 , 8),
			to_signed( -19 , 8),
			to_signed( -6 , 8),
			to_signed( -13 , 8),
			to_signed( -19 , 8),
			to_signed( -16 , 8),
			to_signed( 29 , 8),
			to_signed( -2 , 8),
			to_signed( -4 , 8),
			to_signed( -12 , 8),
			to_signed( 16 , 8),
			to_signed( 14 , 8),
			to_signed( 9 , 8),
			to_signed( -1 , 8),
			to_signed( -22 , 8),
			to_signed( -3 , 8),
			to_signed( 7 , 8),
			to_signed( 7 , 8),
			to_signed( -15 , 8),
			to_signed( 10 , 8),
			to_signed( 26 , 8),
			to_signed( 21 , 8),
			to_signed( -10 , 8),
			to_signed( -32 , 8),
			to_signed( -31 , 8),
			to_signed( 35 , 8),
			to_signed( 0 , 8),
			to_signed( -1 , 8),
			to_signed( 18 , 8),
			to_signed( 26 , 8),
			to_signed( 41 , 8),
			to_signed( -8 , 8),
			to_signed( -16 , 8),
			to_signed( -1 , 8),
			to_signed( -9 , 8),
			to_signed( 8 , 8),
			to_signed( -16 , 8),
			to_signed( -10 , 8),
			to_signed( 3 , 8),
			to_signed( 13 , 8),
			to_signed( -2 , 8),
			to_signed( -33 , 8),
			to_signed( -3 , 8),
			to_signed( 16 , 8),
			to_signed( 46 , 8),
			to_signed( 22 , 8),
			to_signed( 3 , 8),
			to_signed( 19 , 8),
			to_signed( 33 , 8),
			to_signed( 31 , 8),
			to_signed( 4 , 8),
			to_signed( 6 , 8),
			to_signed( 9 , 8),
			to_signed( 1 , 8),
			to_signed( -1 , 8),
			to_signed( -17 , 8),
			to_signed( 27 , 8),
			to_signed( 34 , 8),
			to_signed( -13 , 8),
			to_signed( -13 , 8),
			to_signed( -34 , 8),
			to_signed( 8 , 8),
			to_signed( 9 , 8),
			to_signed( -2 , 8),
			to_signed( -3 , 8),
			to_signed( -2 , 8),
			to_signed( 7 , 8),
			to_signed( 15 , 8),
			to_signed( 13 , 8),
			to_signed( 15 , 8),
			to_signed( 20 , 8),
			to_signed( -34 , 8),
			to_signed( 3 , 8),
			to_signed( -26 , 8),
			to_signed( -10 , 8),
			to_signed( -12 , 8),
			to_signed( -22 , 8),
			to_signed( 8 , 8),
			to_signed( -5 , 8),
			to_signed( 5 , 8),
			to_signed( 0 , 8),
			to_signed( -26 , 8),
			to_signed( 31 , 8),
			to_signed( 14 , 8),
			to_signed( 7 , 8),
			to_signed( -3 , 8),
			to_signed( -13 , 8),
			to_signed( 10 , 8),
			to_signed( 44 , 8),
			to_signed( 34 , 8),
			to_signed( 10 , 8),
			to_signed( -55 , 8),
			to_signed( 12 , 8),
			to_signed( 38 , 8),
			to_signed( 60 , 8),
			to_signed( 16 , 8),
			to_signed( -29 , 8),
			to_signed( 5 , 8),
			to_signed( 17 , 8),
			to_signed( 49 , 8),
			to_signed( 9 , 8),
			to_signed( 21 , 8),
			to_signed( 15 , 8),
			to_signed( 22 , 8),
			to_signed( 16 , 8),
			to_signed( 13 , 8),
			to_signed( -4 , 8),
			to_signed( -1 , 8),
			to_signed( -1 , 8),
			to_signed( 4 , 8),
			to_signed( -4 , 8),
			to_signed( -5 , 8),
			to_signed( 3 , 8),
			to_signed( -1 , 8),
			to_signed( -7 , 8),
			to_signed( -4 , 8),
			to_signed( -1 , 8),
			to_signed( -1 , 8),
			to_signed( -2 , 8),
			to_signed( -5 , 8),
			to_signed( -1 , 8),
			to_signed( -5 , 8),
			to_signed( 9 , 8),
			to_signed( 1 , 8),
			to_signed( 4 , 8),
			to_signed( 7 , 8),
			to_signed( -3 , 8),
			to_signed( -4 , 8),
			to_signed( 4 , 8),
			to_signed( -4 , 8),
			to_signed( 0 , 8),
			to_signed( 16 , 8),
			to_signed( 9 , 8),
			to_signed( -9 , 8),
			to_signed( 4 , 8),
			to_signed( -15 , 8),
			to_signed( 7 , 8),
			to_signed( -3 , 8),
			to_signed( -8 , 8),
			to_signed( -15 , 8),
			to_signed( 0 , 8),
			to_signed( -1 , 8),
			to_signed( -6 , 8),
			to_signed( -8 , 8),
			to_signed( 23 , 8),
			to_signed( 30 , 8),
			to_signed( -29 , 8),
			to_signed( -30 , 8),
			to_signed( 12 , 8),
			to_signed( -1 , 8),
			to_signed( 8 , 8),
			to_signed( -10 , 8),
			to_signed( 10 , 8),
			to_signed( -12 , 8),
			to_signed( -24 , 8),
			to_signed( -16 , 8),
			to_signed( 23 , 8),
			to_signed( 16 , 8),
			to_signed( 19 , 8),
			to_signed( -8 , 8),
			to_signed( 1 , 8),
			to_signed( 8 , 8),
			to_signed( 2 , 8),
			to_signed( 27 , 8),
			to_signed( 5 , 8),
			to_signed( -11 , 8),
			to_signed( 12 , 8),
			to_signed( 7 , 8),
			to_signed( -15 , 8),
			to_signed( 25 , 8),
			to_signed( 37 , 8),
			to_signed( -6 , 8),
			to_signed( -34 , 8),
			to_signed( -50 , 8),
			to_signed( -14 , 8),
			to_signed( -14 , 8),
			to_signed( -9 , 8),
			to_signed( -39 , 8),
			to_signed( 14 , 8),
			to_signed( -11 , 8),
			to_signed( -35 , 8),
			to_signed( 14 , 8),
			to_signed( 30 , 8),
			to_signed( 39 , 8),
			to_signed( 50 , 8),
			to_signed( 50 , 8),
			to_signed( -34 , 8),
			to_signed( -39 , 8),
			to_signed( -14 , 8),
			to_signed( 4 , 8),
			to_signed( 7 , 8),
			to_signed( 0 , 8),
			to_signed( -16 , 8),
			to_signed( -9 , 8),
			to_signed( 6 , 8),
			to_signed( 1 , 8),
			to_signed( 13 , 8),
			to_signed( -1 , 8),
			to_signed( 3 , 8),
			to_signed( -17 , 8),
			to_signed( -15 , 8),
			to_signed( -14 , 8),
			to_signed( -3 , 8),
			to_signed( -13 , 8),
			to_signed( 5 , 8),
			to_signed( -6 , 8),
			to_signed( 4 , 8),
			to_signed( -24 , 8),
			to_signed( 8 , 8),
			to_signed( -16 , 8),
			to_signed( -6 , 8),
			to_signed( 21 , 8),
			to_signed( -10 , 8),
			to_signed( -3 , 8),
			to_signed( -5 , 8),
			to_signed( 4 , 8),
			to_signed( 13 , 8),
			to_signed( 4 , 8),
			to_signed( -14 , 8),
			to_signed( -20 , 8),
			to_signed( 14 , 8),
			to_signed( 6 , 8),
			to_signed( 11 , 8),
			to_signed( 15 , 8),
			to_signed( 2 , 8),
			to_signed( -4 , 8),
			to_signed( -5 , 8),
			to_signed( -41 , 8),
			to_signed( -30 , 8),
			to_signed( -29 , 8),
			to_signed( -27 , 8),
			to_signed( -4 , 8),
			to_signed( -18 , 8),
			to_signed( -30 , 8),
			to_signed( -45 , 8),
			to_signed( -44 , 8),
			to_signed( -2 , 8),
			to_signed( 13 , 8),
			to_signed( 1 , 8),
			to_signed( 10 , 8),
			to_signed( -18 , 8),
			to_signed( -7 , 8),
			to_signed( 21 , 8),
			to_signed( 16 , 8),
			to_signed( 0 , 8),
			to_signed( 15 , 8),
			to_signed( 7 , 8),
			to_signed( 22 , 8),
			to_signed( 8 , 8),
			to_signed( 8 , 8),
			to_signed( 4 , 8),
			to_signed( 4 , 8),
			to_signed( 1 , 8),
			to_signed( 9 , 8),
			to_signed( -10 , 8),
			to_signed( -8 , 8)
	);
	signal weight : signed(7 downto 0);
	signal datas  : data_array(0 to 399) := (
			to_unsigned( 17 , 8),
			to_unsigned( 31 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 21 , 8),
			to_unsigned( 14 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 42 , 8),
			to_unsigned( 59 , 8),
			to_unsigned( 51 , 8),
			to_unsigned( 12 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 63 , 8),
			to_unsigned( 76 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 17 , 8),
			to_unsigned( 44 , 8),
			to_unsigned( 73 , 8),
			to_unsigned( 26 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 12 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 19 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 7 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 23 , 8),
			to_unsigned( 28 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 18 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 36 , 8),
			to_unsigned( 40 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 29 , 8),
			to_unsigned( 11 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 22 , 8),
			to_unsigned( 13 , 8),
			to_unsigned( 1 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 19 , 8),
			to_unsigned( 19 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 56 , 8),
			to_unsigned( 53 , 8),
			to_unsigned( 44 , 8),
			to_unsigned( 54 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 22 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 31 , 8),
			to_unsigned( 51 , 8),
			to_unsigned( 31 , 8),
			to_unsigned( 23 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 18 , 8),
			to_unsigned( 42 , 8),
			to_unsigned( 18 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 40 , 8),
			to_unsigned( 30 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 38 , 8),
			to_unsigned( 26 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 35 , 8),
			to_unsigned( 31 , 8),
			to_unsigned( 41 , 8),
			to_unsigned( 68 , 8),
			to_unsigned( 37 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 19 , 8),
			to_unsigned( 38 , 8),
			to_unsigned( 14 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 30 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 20 , 8),
			to_unsigned( 14 , 8),
			to_unsigned( 13 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 20 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 5 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 7 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 20 , 8),
			to_unsigned( 21 , 8),
			to_unsigned( 17 , 8),
			to_unsigned( 23 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 25 , 8),
			to_unsigned( 33 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 64 , 8),
			to_unsigned( 54 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 72 , 8),
			to_unsigned( 49 , 8),
			to_unsigned( 1 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 48 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 80 , 8),
			to_unsigned( 115 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 44 , 8),
			to_unsigned( 121 , 8),
			to_unsigned( 86 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 120 , 8),
			to_unsigned( 127 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 23 , 8),
			to_unsigned( 106 , 8),
			to_unsigned( 55 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 22 , 8),
			to_unsigned( 41 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 5 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 43 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 5 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 50 , 8),
			to_unsigned( 54 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 18 , 8),
			to_unsigned( 9 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 11 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 4 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 26 , 8),
			to_unsigned( 24 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 8 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 28 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 45 , 8),
			to_unsigned( 37 , 8),
			to_unsigned( 54 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 25 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 26 , 8),
			to_unsigned( 31 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 5 , 8),
			to_unsigned( 9 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 20 , 8),
			to_unsigned( 2 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 24 , 8),
			to_unsigned( 10 , 8),
			to_unsigned( 12 , 8),
			to_unsigned( 23 , 8),
			to_unsigned( 32 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 35 , 8),
			to_unsigned( 30 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 7 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 16 , 8),
			to_unsigned( 36 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 21 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 1 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 15 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 13 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 3 , 8),
			to_unsigned( 25 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 22 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 22 , 8),
			to_unsigned( 7 , 8),
			to_unsigned( 33 , 8),
			to_unsigned( 86 , 8),
			to_unsigned( 1 , 8),
			to_unsigned( 9 , 8),
			to_unsigned( 6 , 8),
			to_unsigned( 75 , 8),
			to_unsigned( 104 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 61 , 8),
			to_unsigned( 53 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 38 , 8),
			to_unsigned( 58 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 34 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8),
			to_unsigned( 0 , 8)
	);
	signal data : unsigned(7 downto 0);
	signal bias : signed(31 downto 0) := to_signed(97, 32);

	constant scale : integer := integer(0.0023508628364652395 * 2**16); -- Scale value in fixed-point (scaled by 256)

	signal index : integer := 0;

begin

		U1 : channel_layer_5 port map(
			clka           => clka,
			resetn         => resetn,
			start          => start,
			finish         => finish,
			weight         => weight,
			bias           => bias,
			data           => data,
			compute_output => compute_output,
			scale          => scale
		);

	clka_process : process
	begin
		while true loop
			clka <= '0';
			wait for CLK_PERIOD / 2;
			clka <= '1';
			wait for CLK_PERIOD / 2;
		end loop;
	end process;

	resetn_process : process(clka)
	begin
		if rising_edge(clka) then
			if resetn_flag = 0 then
				resetn      <= '0';
				resetn_flag <= 1;
			else
				resetn <= '1';
			end if;
		end if;
	end process;

	start_process : process(clka)
	begin
		if rising_edge(clka) and resetn = '1' then
			if finish = '1' then
				start_flag <= 0;
			elsif start_flag = 0 then
				if index < 400 then
					weight <= weights(index);
					data   <= datas(index);
					index  <= index + 1;
				end if;

				start      <= '1';
				start_flag <= 1;
			else
				start <= '0';
			end if;
		end if;
	end process;

	--	main_process : process(clka)
	--	begin
	--		if resetn = '1' then
	--			if rising_edge(clka) then
	--				if finish = '1' then

	--				end if;

--			end if;
--		end if;
--	end process;
end Behavioral;